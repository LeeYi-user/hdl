LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY N_COUNTER is
	PORT( CLK: IN STD_LOGIC;
			Q: OUT STD_LOGIC);
END N_COUNTER;

ARCHITECTURE a OF N_COUNTER IS
	SIGNAL QN : STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL RESET:STD_LOGIC;
BEGIN
	PROCESS (CLK)
		BEGIN
			IF RESET='1' THEN QN<="0000";
			ELSIF CLK'event AND CLK='1' THEN QN <= QN+1;
			END IF;
	END PROCESS;
	RESET<='1' WHEN QN=10 ELSE '0';
	Q<=QN(3);
END a;
